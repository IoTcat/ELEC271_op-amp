* C:\Users\ushio\OneDrive\study\uol\ELEC271\ex5\part1\part1.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 05 17:50:20 2020



** Analysis setup **
.DC LIN V_Vce 0V 20V 0.5V 
+ LIN I_Ib 0A 40e-6A 4e-6A 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "part1.net"
.INC "part1.als"


.probe


.END
